--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:13:28 08/28/2018
-- Design Name:   
-- Module Name:   /home/sd/Desktop/Trabalho1SD_ULA/testSomadorDe1bitDaRapeize.vhd
-- Project Name:  Trabalho1SD_ULA
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: fullAdder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY testFullAdder IS
END testFullAdder;
 
ARCHITECTURE behavior OF testFullAdder IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT fullAdder
    PORT(
         a : IN  std_logic;
         b : IN  std_logic;
         carryIn : IN  std_logic;
         s : OUT  std_logic;
         carryOut : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic := '0';
   signal b : std_logic := '0';
   signal carryIn : std_logic := '0';

 	--Outputs
   signal s : std_logic;
   signal carryOut : std_logic;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: fullAdder PORT MAP (
          a => a,
          b => b,
          carryIn => carryIn,
          s => s,
          carryOut => carryOut
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

    --  wait for <clock>_period*10;

      -- insert stimulus here 
		
		a <= '0';
		b <= '0';
		carryIn <= '0';
		wait for 10 ns;

		a <= '0';
		b <= '0';
		carryIn <= '1';
		wait for 10 ns;

		a <= '0';
		b <= '1';
		carryIn <= '0';
		wait for 10 ns;
		
		a <= '0';
		b <= '1';
		carryIn <= '1';
		wait for 10 ns;
		
		a <= '1';
		b <= '0';
		carryIn <= '0';
		wait for 10 ns;
		
		a <= '1';
		b <= '0';
		carryIn <= '1';
		wait for 10 ns;
		
		a <= '1';
		b <= '1';
		carryIn <= '0';
		wait for 10 ns;
		
		a <= '1';
		b <= '1';
		carryIn <= '1';
		wait for 10 ns;
      wait;
   end process;

END;
